/* 
wreg_dst_sel控制将被写入的寄存器的编号的来源，
	0来自Instr[20:16](Rt)，1来自Instr[15:11](Rd)
wrbck_sel控制将被写入的寄存器的数据的来源
	0来自aluout，1来自内存输出
*/
module multicyc_mcu (
	input logic clk, reset, 
	input logic [5:0] opcode,

	output logic mem_addr_sel, ir_we,
	output logic alu_srca_sel, 
	output logic [1:0]alu_srcb_sel, 
	output logic [1:0] aluop, 
	output logic mem_rd, mem_wr, 
	reg_we, pc_we, 
	wreg_dst_sel, wrbck_data_sel
);

import ALUops::*;
import Opcodes::*;
import MultcycCtrl::*;



logic [3:0] curr_state;
logic [3:0] next_state;

always_ff @( posedge clk ) begin
	if (reset) curr_state <= 4'b0000;
	else 	   curr_state <= next_state;
end

always_comb begin 
	{mem_addr_sel, ir_we} = 2'b0;
	{alu_srca_sel, alu_srcb_sel, aluop} = 5'b0;
	{mem_rd, mem_wr, reg_we, pc_we, wreg_dst_sel, wrbck_data_sel} = 6'b0;

	case (curr_state)
		Fetch: begin
			next_state = Decode;
			mem_addr_sel = AddrPC;
			alu_srca_sel = SrcaPC;
			alu_srcb_sel = Four;
			aluop = ALUop_ADD;
			ir_we = 1;
			pc_we = 1;	end
		Decode: begin
			if (opcode == LW || opcode == SW) next_state = MemAddr;
			else if (opcode == RR) next_state = RRExec;
			else if (opcode == ADDI) next_state = AddiExec;
			else if (opcode == ADDIU) next_state = AddiuExec;
			else next_state = 0; end
		MemAddr: begin
			next_state = opcode == LW ? MemRd : MemWr;
			alu_srca_sel = SrcaRs;
			alu_srcb_sel = SrcbImm;
			aluop = ALUop_ADD; end
		MemRd: begin
			next_state = MemWrbck;
			mem_addr_sel = AddrALUout;
		end
		MemWr: begin
			next_state = Fetch;
			mem_addr_sel = AddrALUout;
			mem_wr = 1; end
		MemWrbck: begin
			next_state = Fetch;
			wreg_dst_sel = WrRt;
			wrbck_data_sel = MemData;
			reg_we = 1; end
		RRExec: begin
			next_state = ALURRWrbck;
			alu_srca_sel = SrcaRs;
			alu_srcb_sel = SrcbRt;
			aluop = ALUop_RR; end
		ALURRWrbck: begin
			next_state = Fetch;
			wreg_dst_sel = WrRd;
			wrbck_data_sel = ALUout;
			reg_we = 1; end
		AddiExec: begin
			next_state = ALURIWrbck;
			alu_srca_sel = SrcaRs;
			alu_srcb_sel = SrcbImm;
			aluop = ALUop_ADD; end
		AddiuExec: begin
			next_state = ALURIWrbck;
			alu_srca_sel = SrcaRs;
			alu_srcb_sel = SrcbImm;
			aluop = ALUop_ADDU; end
		ALURIWrbck: begin
			next_state = Fetch;
			wreg_dst_sel = WrRt;
			wrbck_data_sel = ALUout;
			reg_we = 1;
		end
			
		default: ;
	endcase
end
	
endmodule
